module scr1_tb_log_cmd();

always_ff @(posedge scr1_top_tb_ahb.i_top.i_imem_ahb.clk) begin
    if (scr1_top_tb_ahb.i_top.i_imem_ahb.imem_resp == 2'b01) begin
        // valid data from ahb router
        if (
            (scr1_top_tb_ahb.i_top.i_imem_ahb.imem_rdata[31 : 0] == 32'h1DD19963)
        ) begin
            // detect and command
            $display("PC: %04h",scr1_top_tb_ahb.i_top.i_core_top.i_pipe_top.curr_pc);
        end
    end
end

endmodule